`timescale 1us/1us

module dff (
  input logic clk, d,
  output logic q
);

// Internal logic

endmodule
